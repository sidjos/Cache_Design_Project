-- Level 1 Cache
