library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.eecs361_gates.all;
use work.eecs361.all;

entity main_memory is
	generic ( mem_file: string);
	port (
		clk:     		in std_logic; 
		reset:		in std_logic; 
		address:		in std_logic_vector(31 downto 0); 
		L2_Miss: 	in std_logic;
		main_write: 	in std_logic;
		data_in: 	in std_logic_vector (31 downto 0);
		data_valid: 	out std_logic;
		data_out_with_tag: 	out std_logic_vector(2069 downto 0)
	);
end main_memory;

architecture structural of main_memory is

signal mux0,mux1,mux2,mux3,mux4,shifter,fulladder1, data_out_sig: std_logic_vector(2047 downto 0);
signal mux6: std_logic_vector(9 downto 0);
signal syncram0,counter,pc0,counter_minus_one,fulladder2: std_logic_vector(31 downto 0);
signal not0,and0,counter_minus_one_to_be_64,clk_with_stop,clk_with_stop_and_trigger,not_clk_with_stop_and_trigger: std_logic;


begin
        
   

   --valid 
   data_valid <= counter_minus_one_to_be_64;
   and0_map: and_gate port map (x=>counter_minus_one(6), y=>counter_minus_one(0), z=>counter_minus_one_to_be_64);
   or0_map:  or_gate port map (x=>clk, y=>counter_minus_one_to_be_64, z=>clk_with_stop);
   and1_map:  or_gate port map (x=>clk_with_stop, y=>L2_Miss, z=>clk_with_stop_and_trigger);
   not0_map:	not_gate port map (x=>clk_with_stop_and_trigger,z=>not_clk_with_stop_and_trigger);


   --main memory 
   mux6_map: 	mux_n generic map (n=>10) port map (sel=>main_write, src0=>B"0000000000", src1=>address(9 downto 0), z=>mux6);

   syncram_map:	syncram generic map (mem_file => mem_file)
				port map (clk=>clk_with_stop_and_trigger, cs=>'1', oe=>'1', we=>main_write, addr(31 downto 10)=>address(31 downto 10), addr(9 downto 0)=>mux6, din=>data_in, dout=>syncram0);
  
   --32 bits counter (positive edge)
   fulladder0_map:  fulladder_32 port map (cin=>'0', x=>pc0, y=>B"00000000000000000000000000000001", z=>counter);
   generate_memory0: for i in 0 to 31 generate
   map_memory_reg0: dffr_a port map (clk=>clk_with_stop_and_trigger, arst=>reset, aload=>'0', adata=>'0', d=>counter(i), enable=>'1',q=>pc0(i));
   end generate generate_memory0;
   
    fulladder2_map:  fulladder_32 port map (cin=>'0', x=>pc0, y=>B"11111111111111111111111111111111", z=>counter_minus_one);
   --temporary 256 bytes Registers (negative edge)
   --1024-bit
   mux0_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(5), 
   							   src0(31 downto 0)=>syncram0,
   							   src0(2047 downto 32)=>B"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
   							   src1(1055 downto 1024)=>syncram0,
   							   src1(2047 downto 1056)=>B"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
   							   src1(511 downto 0)=>B"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
   							   src1(1023 downto 512)=>B"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
   							   z=>mux0);
   --512-bit
   mux1_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(4), src0=>mux0, src1(2047 downto 512)=>mux0(1535 downto 0),src1(511 downto 0)=>B"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", z=>mux1);
   --256-bit
   mux2_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(3), src0=>mux1, src1(2047 downto 256)=>mux1(1791 downto 0),src1(255 downto 0)=>B"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", z=>mux2);
   --128-bit
   mux3_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(2), src0=>mux2, src1(2047 downto 128)=>mux2(1919 downto 0),src1(127 downto 0)=>B"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", z=>mux3);
   --64-bit
   mux4_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(1), src0=>mux3, src1(2047 downto 64)=>mux3(1983 downto 0),src1(63 downto 0)=>B"0000000000000000000000000000000000000000000000000000000000000000", z=>mux4);
   --32-bit
   mux5_map:	mux_n generic map (n=>2048)	 port map (sel=>counter_minus_one(0), src0=>mux4, src1(2047 downto 32)=>mux4(2015 downto 0),src1(31 downto 0)=>B"00000000000000000000000000000000", z=>shifter);
   
   data_out_with_tag <= address(31 downto 10) & data_out_sig;
   
   fulladder1_map:  fulladder_n generic map (n=>2048) port map (cin=>'0', x=>data_out_sig, y=>shifter, z=>fulladder1);

   generate_memory1: for i in 0 to 2047 generate
   map_memory_reg1: dffr_a port map (clk=>not_clk_with_stop_and_trigger, arst=>reset,aload=>'0', adata=>'0', d=>fulladder1(i), enable=>'1',q=>data_out_sig(i));
   end generate generate_memory1;
   
end architecture structural;

